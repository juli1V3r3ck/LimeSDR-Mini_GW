// factory.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module factory (
		input  wire [20:0] bridge_0_address,     // bridge_0.address
		input  wire [3:0]  bridge_0_byte_enable, //         .byte_enable
		input  wire        bridge_0_read,        //         .read
		input  wire        bridge_0_write,       //         .write
		input  wire [31:0] bridge_0_write_data,  //         .write_data
		output wire        bridge_0_acknowledge, //         .acknowledge
		output wire [31:0] bridge_0_read_data,   //         .read_data
		input  wire        clk_clk,              //      clk.clk
		output wire [31:0] extfifo_of_d,         //  extfifo.of_d
		output wire        extfifo_of_wr,        //         .of_wr
		input  wire        extfifo_of_wrfull,    //         .of_wrfull
		input  wire [31:0] extfifo_if_d,         //         .if_d
		output wire        extfifo_if_rd,        //         .if_rd
		input  wire        extfifo_if_rdempty,   //         .if_rdempty
		output wire        extfifo_fifo_rst,     //         .fifo_rst
		output wire [7:0]  pio_0_export,         //    pio_0.export
		input  wire        reset_reset_n,        //    reset.reset_n
		inout  wire        scl_export,           //      scl.export
		inout  wire        sda_export            //      sda.export
	);

	wire  [31:0] bridge_0_avalon_master_readdata;                              // mm_interconnect_0:bridge_0_avalon_master_readdata -> bridge_0:avalon_readdata
	wire         bridge_0_avalon_master_waitrequest;                           // mm_interconnect_0:bridge_0_avalon_master_waitrequest -> bridge_0:avalon_waitrequest
	wire   [3:0] bridge_0_avalon_master_byteenable;                            // bridge_0:avalon_byteenable -> mm_interconnect_0:bridge_0_avalon_master_byteenable
	wire         bridge_0_avalon_master_read;                                  // bridge_0:avalon_read -> mm_interconnect_0:bridge_0_avalon_master_read
	wire  [20:0] bridge_0_avalon_master_address;                               // bridge_0:avalon_address -> mm_interconnect_0:bridge_0_avalon_master_address
	wire         bridge_0_avalon_master_write;                                 // bridge_0:avalon_write -> mm_interconnect_0:bridge_0_avalon_master_write
	wire  [31:0] bridge_0_avalon_master_writedata;                             // bridge_0:avalon_writedata -> mm_interconnect_0:bridge_0_avalon_master_writedata
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_readdata;                // dual_boot_0:avmm_rcv_readdata -> mm_interconnect_0:dual_boot_0_avalon_readdata
	wire   [2:0] mm_interconnect_0_dual_boot_0_avalon_address;                 // mm_interconnect_0:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	wire         mm_interconnect_0_dual_boot_0_avalon_read;                    // mm_interconnect_0:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	wire         mm_interconnect_0_dual_boot_0_avalon_write;                   // mm_interconnect_0:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_0_dual_boot_0_avalon_writedata;               // mm_interconnect_0:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect;  // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata;    // i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest; // i2c_opencores_0:wb_ack_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address;     // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write;       // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata;   // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata;             // avs_fifo_int_0:avs_s0_readdata -> mm_interconnect_0:avs_fifo_int_0_avs_s0_readdata
	wire         mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest;          // avs_fifo_int_0:avs_s0_waitrequest -> mm_interconnect_0:avs_fifo_int_0_avs_s0_waitrequest
	wire   [7:0] mm_interconnect_0_avs_fifo_int_0_avs_s0_address;              // mm_interconnect_0:avs_fifo_int_0_avs_s0_address -> avs_fifo_int_0:avs_s0_address
	wire         mm_interconnect_0_avs_fifo_int_0_avs_s0_read;                 // mm_interconnect_0:avs_fifo_int_0_avs_s0_read -> avs_fifo_int_0:avs_s0_read
	wire         mm_interconnect_0_avs_fifo_int_0_avs_s0_write;                // mm_interconnect_0:avs_fifo_int_0_avs_s0_write -> avs_fifo_int_0:avs_s0_write
	wire  [31:0] mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata;            // mm_interconnect_0:avs_fifo_int_0_avs_s0_writedata -> avs_fifo_int_0:avs_s0_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                 // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                    // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                   // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;               // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;               // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;            // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [17:0] mm_interconnect_0_onchip_flash_0_data_address;                // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                   // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;          // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                  // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;              // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;             // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire         mm_interconnect_0_pio_0_s1_chipselect;                        // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                          // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_0_s1_address;                           // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                             // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                         // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [avs_fifo_int_0:reset_reset, bridge_0:reset, dual_boot_0:nreset, i2c_opencores_0:wb_rst_i, mm_interconnect_0:bridge_0_reset_reset_bridge_in_reset_reset, onchip_flash_0:reset_n, pio_0:reset_n]

	avs_fifo_int avs_fifo_int_0 (
		.avs_s0_address     (mm_interconnect_0_avs_fifo_int_0_avs_s0_address),     // avs_s0.address
		.avs_s0_read        (mm_interconnect_0_avs_fifo_int_0_avs_s0_read),        //       .read
		.avs_s0_readdata    (mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata),    //       .readdata
		.avs_s0_write       (mm_interconnect_0_avs_fifo_int_0_avs_s0_write),       //       .write
		.avs_s0_writedata   (mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata),   //       .writedata
		.avs_s0_waitrequest (mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest), //       .waitrequest
		.clock_clk          (clk_clk),                                             //  clock.clk
		.reset_reset        (rst_controller_reset_out_reset),                      //  reset.reset
		.of_d               (extfifo_of_d),                                        //    coe.of_d
		.of_wr              (extfifo_of_wr),                                       //       .of_wr
		.of_wrfull          (extfifo_of_wrfull),                                   //       .of_wrfull
		.if_d               (extfifo_if_d),                                        //       .if_d
		.if_rd              (extfifo_if_rd),                                       //       .if_rd
		.if_rdempty         (extfifo_if_rdempty),                                  //       .if_rdempty
		.fifo_rst           (extfifo_fifo_rst)                                     //       .fifo_rst
	);

	factory_bridge_0 bridge_0 (
		.clk                (clk_clk),                            //                clk.clk
		.reset              (rst_controller_reset_out_reset),     //              reset.reset
		.avalon_readdata    (bridge_0_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_0_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_0_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_0_avalon_master_read),        //                   .read
		.avalon_write       (bridge_0_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_0_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_0_avalon_master_address),     //                   .address
		.address            (bridge_0_address),                   // external_interface.export
		.byte_enable        (bridge_0_byte_enable),               //                   .export
		.read               (bridge_0_read),                      //                   .export
		.write              (bridge_0_write),                     //                   .export
		.write_data         (bridge_0_write_data),                //                   .export
		.acknowledge        (bridge_0_acknowledge),               //                   .export
		.read_data          (bridge_0_read_data)                  //                   .export
	);

	altera_dual_boot #(
		.INTENDED_DEVICE_FAMILY ("MAX 10"),
		.CONFIG_CYCLE           (15),
		.RESET_TIMER_CYCLE      (21)
	) dual_boot_0 (
		.clk                (clk_clk),                                        //    clk.clk
		.nreset             (~rst_controller_reset_out_reset),                // nreset.reset_n
		.avmm_rcv_address   (mm_interconnect_0_dual_boot_0_avalon_address),   // avalon.address
		.avmm_rcv_read      (mm_interconnect_0_dual_boot_0_avalon_read),      //       .read
		.avmm_rcv_writedata (mm_interconnect_0_dual_boot_0_avalon_writedata), //       .writedata
		.avmm_rcv_write     (mm_interconnect_0_dual_boot_0_avalon_write),     //       .write
		.avmm_rcv_readdata  (mm_interconnect_0_dual_boot_0_avalon_readdata)   //       .readdata
	);

	i2c_opencores i2c_opencores_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (scl_export),                                                   //       export_scl.export
		.sda_pad_io (sda_export),                                                   //       export_sda.export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  ()                                                              // interrupt_sender.irq
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M16SAU169I7G"),
		.DEVICE_ID                           ("16"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (47103),
		.SECTOR4_START_ADDR                  (47104),
		.SECTOR4_END_ADDR                    (75775),
		.SECTOR5_START_ADDR                  (75776),
		.SECTOR5_END_ADDR                    (143359),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (143359),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (8191),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (143359),
		.ADDR_RANGE2_END_ADDR                (143359),
		.ADDR_RANGE1_OFFSET                  (1024),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (18),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (10),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (48),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (14000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (12200),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("True"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) onchip_flash_0 (
		.clock                   (clk_clk),                                             //    clk.clk
		.reset_n                 (~rst_controller_reset_out_reset),                     // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	factory_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_export)                           // external_connection.export
	);

	factory_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                              (clk_clk),                                                       //                            clk_0_clk.clk
		.bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // bridge_0_reset_reset_bridge_in_reset.reset
		.bridge_0_avalon_master_address             (bridge_0_avalon_master_address),                                //               bridge_0_avalon_master.address
		.bridge_0_avalon_master_waitrequest         (bridge_0_avalon_master_waitrequest),                            //                                     .waitrequest
		.bridge_0_avalon_master_byteenable          (bridge_0_avalon_master_byteenable),                             //                                     .byteenable
		.bridge_0_avalon_master_read                (bridge_0_avalon_master_read),                                   //                                     .read
		.bridge_0_avalon_master_readdata            (bridge_0_avalon_master_readdata),                               //                                     .readdata
		.bridge_0_avalon_master_write               (bridge_0_avalon_master_write),                                  //                                     .write
		.bridge_0_avalon_master_writedata           (bridge_0_avalon_master_writedata),                              //                                     .writedata
		.avs_fifo_int_0_avs_s0_address              (mm_interconnect_0_avs_fifo_int_0_avs_s0_address),               //                avs_fifo_int_0_avs_s0.address
		.avs_fifo_int_0_avs_s0_write                (mm_interconnect_0_avs_fifo_int_0_avs_s0_write),                 //                                     .write
		.avs_fifo_int_0_avs_s0_read                 (mm_interconnect_0_avs_fifo_int_0_avs_s0_read),                  //                                     .read
		.avs_fifo_int_0_avs_s0_readdata             (mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata),              //                                     .readdata
		.avs_fifo_int_0_avs_s0_writedata            (mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata),             //                                     .writedata
		.avs_fifo_int_0_avs_s0_waitrequest          (mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest),           //                                     .waitrequest
		.dual_boot_0_avalon_address                 (mm_interconnect_0_dual_boot_0_avalon_address),                  //                   dual_boot_0_avalon.address
		.dual_boot_0_avalon_write                   (mm_interconnect_0_dual_boot_0_avalon_write),                    //                                     .write
		.dual_boot_0_avalon_read                    (mm_interconnect_0_dual_boot_0_avalon_read),                     //                                     .read
		.dual_boot_0_avalon_readdata                (mm_interconnect_0_dual_boot_0_avalon_readdata),                 //                                     .readdata
		.dual_boot_0_avalon_writedata               (mm_interconnect_0_dual_boot_0_avalon_writedata),                //                                     .writedata
		.i2c_opencores_0_avalon_slave_0_address     (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),      //       i2c_opencores_0_avalon_slave_0.address
		.i2c_opencores_0_avalon_slave_0_write       (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),        //                                     .write
		.i2c_opencores_0_avalon_slave_0_readdata    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),     //                                     .readdata
		.i2c_opencores_0_avalon_slave_0_writedata   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),    //                                     .writedata
		.i2c_opencores_0_avalon_slave_0_waitrequest (~mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                                     .waitrequest
		.i2c_opencores_0_avalon_slave_0_chipselect  (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),   //                                     .chipselect
		.onchip_flash_0_csr_address                 (mm_interconnect_0_onchip_flash_0_csr_address),                  //                   onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                   (mm_interconnect_0_onchip_flash_0_csr_write),                    //                                     .write
		.onchip_flash_0_csr_read                    (mm_interconnect_0_onchip_flash_0_csr_read),                     //                                     .read
		.onchip_flash_0_csr_readdata                (mm_interconnect_0_onchip_flash_0_csr_readdata),                 //                                     .readdata
		.onchip_flash_0_csr_writedata               (mm_interconnect_0_onchip_flash_0_csr_writedata),                //                                     .writedata
		.onchip_flash_0_data_address                (mm_interconnect_0_onchip_flash_0_data_address),                 //                  onchip_flash_0_data.address
		.onchip_flash_0_data_write                  (mm_interconnect_0_onchip_flash_0_data_write),                   //                                     .write
		.onchip_flash_0_data_read                   (mm_interconnect_0_onchip_flash_0_data_read),                    //                                     .read
		.onchip_flash_0_data_readdata               (mm_interconnect_0_onchip_flash_0_data_readdata),                //                                     .readdata
		.onchip_flash_0_data_writedata              (mm_interconnect_0_onchip_flash_0_data_writedata),               //                                     .writedata
		.onchip_flash_0_data_burstcount             (mm_interconnect_0_onchip_flash_0_data_burstcount),              //                                     .burstcount
		.onchip_flash_0_data_readdatavalid          (mm_interconnect_0_onchip_flash_0_data_readdatavalid),           //                                     .readdatavalid
		.onchip_flash_0_data_waitrequest            (mm_interconnect_0_onchip_flash_0_data_waitrequest),             //                                     .waitrequest
		.pio_0_s1_address                           (mm_interconnect_0_pio_0_s1_address),                            //                             pio_0_s1.address
		.pio_0_s1_write                             (mm_interconnect_0_pio_0_s1_write),                              //                                     .write
		.pio_0_s1_readdata                          (mm_interconnect_0_pio_0_s1_readdata),                           //                                     .readdata
		.pio_0_s1_writedata                         (mm_interconnect_0_pio_0_s1_writedata),                          //                                     .writedata
		.pio_0_s1_chipselect                        (mm_interconnect_0_pio_0_s1_chipselect)                          //                                     .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
